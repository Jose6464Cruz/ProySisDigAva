----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:05:51 12/08/2019 
-- Design Name: 
-- Module Name:    VGA_DISPLAY - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity VGA_DISPLAY is
   -- Used for the ROM
  Generic
	 ( n : integer := 12;   -- Number of Address bus lines
	   m : integer := 8);   -- Number of Data bus lines
  port (
    Clk : in  STD_LOGIC;
	 Xin : in  STD_LOGIC_VECTOR(9 downto 0); -- Column screen coordinate
	 Yin : in  STD_LOGIC_VECTOR(9 downto 0); -- Row screen coordinate
	 En  : in  STD_LOGIC;                    -- When '1', pixels can be drawn 
	 img : in  STD_LOGIC_VECTOR(2 downto 0);
	 R   : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Red channel
	 G   : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Green channel
	 B   : out STD_LOGIC_VECTOR(1 downto 0));-- 2-bit Blue channel
end VGA_DISPLAY;

architecture Behavioral of VGA_DISPLAY is

  -- Embedded signal to group the colors into 1-byte
  -- The colors will be as follows:
  --  R2 R1 R0 G2 G1 G0 B1 B0
  signal Color :  STD_LOGIC_VECTOR(7 downto 0);
  --signal Address: STD_LOGIC_VECTOR(n-1 downto 0);
  signal Data:    STD_LOGIC_VECTOR(m-1 downto 0);
  signal Address: integer range 0 to (2**n);
  
  -- ROM Declaration
  -- Matrix declaration for ROM
  type type_ROM is array (0 to (2**n) - 1) of STD_LOGIC_VECTOR (m-1 downto 0);
  constant ROM_MOTORCYCLE : type_ROM := 
(x"DC",x"DD",x"00",x"00",x"00",x"DD",x"DC",x"DD",
x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FD",x"DC",x"DC",
x"DC",x"DD",x"FE",x"00",x"FD",x"DC",x"DC",x"DD",
x"00",x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FD",x"DC",x"DC",
x"DD",x"DC",x"FD",x"00",x"FD",x"DC",x"DD",x"DD",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DD",
x"DD",x"DD",x"FE",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"FD",x"DD",x"DD",x"DD",x"FD",x"00",
x"00",x"00",x"DD",x"DD",x"DD",x"DD",x"FE",x"00",
x"00",x"FD",x"DD",x"DD",x"DD",x"DD",x"DD",x"FE",
x"FD",x"DD",x"DD",x"FD",x"00",x"00",x"00",x"FD",
x"DD",x"DD",x"FD",x"00",x"00",x"FD",x"DC",x"DC",
x"00",x"DC",x"FD",x"00",x"DD",x"DC",x"00",x"DC",
x"DD",x"FE",x"DC",x"DC",x"00",x"FE",x"DC",x"DD",
x"FE",x"DD",x"DC",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"FE",x"DC",x"FD",x"FE",x"DC",x"DC",x"FE",
x"00",x"FD",x"DC",x"FE",x"FE",x"FD",x"DC",x"FD",
x"00",x"DD",x"DC",x"DC",x"FE",x"DD",x"DC",x"DC",
x"FD",x"FE",x"DC",x"DD",x"00",x"00",x"DD",x"DC",
x"FD",x"FD",x"DC",x"DD",x"00",x"FE",x"DD",x"DC",
x"00",x"DC",x"FD",x"FE",x"DC",x"FE",x"00",x"DC",
x"DD",x"FE",x"DC",x"FE",x"00",x"DD",x"DC",x"DC",
x"DD",x"DD",x"DC",x"DC",x"00",x"DC",x"DC",x"FD",
x"FE",x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",
x"FE",x"DD",x"DC",x"00",x"00",x"00",x"FE",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"DD",x"DD",x"DC",x"DC",x"FE",x"00",x"DD",x"FE",
x"00",x"DC",x"DC",x"DC",x"DC",x"00",x"00",x"DD",
x"DC",x"DC",x"DC",x"FE",x"00",x"DD",x"DC",x"DC",
x"DD",x"DD",x"DD",x"DD",x"00",x"DC",x"DC",x"FD",
x"FE",x"DC",x"DC",x"00",x"00",x"00",x"00",x"00",
x"FE",x"DC",x"DC",x"00",x"00",x"00",x"FE",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"DD",x"DD",x"DD",x"DD",x"FE",x"00",x"DD",x"00",
x"00",x"FE",x"DC",x"DC",x"DC",x"00",x"00",x"00",
x"DC",x"DC",x"DC",x"FE",x"00",x"DD",x"DC",x"DD",
x"00",x"00",x"FE",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"DD",x"DC",x"00",x"00",x"00",x"FE",x"FE",
x"00",x"DD",x"DC",x"00",x"00",x"00",x"DD",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"00",x"00",x"FE",x"FE",x"00",x"00",x"FE",x"00",
x"00",x"00",x"DC",x"DC",x"FE",x"00",x"00",x"00",
x"DC",x"DC",x"FE",x"00",x"00",x"00",x"DD",x"DC",
x"DD",x"DD",x"DD",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"FE",x"DC",x"DD",x"DD",x"DD",x"DC",x"FE",
x"00",x"FE",x"DC",x"DD",x"DD",x"DD",x"DC",x"FE",
x"00",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"00",x"FE",x"DC",
x"DD",x"DD",x"DC",x"FE",x"00",x"FE",x"DD",x"DD",
x"00",x"00",x"FE",x"FE",x"00",x"00",x"00",x"00",
x"FE",x"FE",x"00",x"00",x"00",x"00",x"00",x"FE",
x"FE",x"FE",x"00",x"00",x"00",x"FE",x"FE",x"FE",
x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",
x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",
x"00",x"FE",x"FE",x"FE",x"00",x"00",x"FE",x"FE",
x"00",x"00",x"FE",x"FE",x"FE",x"00",x"00",x"FE",
x"FE",x"FE",x"FE",x"00",x"00",x"FE",x"FE",x"FE",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DD",x"FE",x"00",x"00",x"FD",x"DC",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FD",x"DC",x"FD",x"00",x"00",x"00",x"00",x"FE",
x"FE",x"00",x"00",x"FE",x"DD",x"DC",x"DC",x"DC",
x"FD",x"00",x"00",x"DD",x"DC",x"DC",x"DC",x"FD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DC",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DD",x"FE",x"FE",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DC",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FE",x"DD",x"DC",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FE",x"DC",x"FD",x"00",x"00",x"00",x"00",x"DD",
x"FE",x"00",x"FE",x"DD",x"DC",x"FE",x"FE",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"DC",x"FD",x"00",x"00",x"DD",x"DC",
x"DC",x"FE",x"FE",x"DC",x"DC",x"FE",x"FE",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FD",x"DC",x"DC",x"DC",x"DC",x"DC",
x"FE",x"00",x"00",x"DD",x"DC",x"DC",x"DC",x"FE",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"DD",x"DD",x"DD",x"DD",x"DD",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DD",
x"DD",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DD",x"FE",x"FE",x"FE",x"DC",x"DC",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"DC",
x"DD",x"00",x"FE",x"DD",x"DD",x"DD",x"DD",x"DD",
x"DD",x"FE",x"00",x"00",x"FE",x"DD",x"DD",x"DD",
x"FE",x"00",x"00",x"00",x"FD",x"DD",x"DD",x"FE",
x"00",x"00",x"00",x"FD",x"DD",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DD",x"00",x"00",x"00",x"DD",x"DC",
x"FE",x"00",x"FE",x"DC",x"DD",x"DD",x"DD",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"DD",x"DD",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"DD",x"DD",x"DC",
x"FE",x"00",x"00",x"FD",x"DD",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"FE",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"FE",x"DD",x"DC",x"00",x"00",x"FE",
x"FE",x"00",x"FD",x"DC",x"DC",x"FE",x"DD",x"DC",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"FE",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"FD",x"DC",x"DC",x"DD",x"DD",x"DD",
x"DD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"FE",x"DD",x"DC",x"00",x"00",x"00",
x"FE",x"00",x"FD",x"DC",x"DC",x"00",x"00",x"FE",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"DD",x"DD",x"DD",
x"DC",x"FE",x"00",x"DD",x"DC",x"DD",x"DD",x"DC",
x"FE",x"00",x"00",x"FD",x"DD",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"FE",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DD",x"00",x"00",x"00",x"DD",
x"DD",x"FE",x"00",x"00",x"FE",x"DD",x"DD",x"DD",
x"FE",x"00",x"00",x"00",x"FD",x"DD",x"DD",x"FE",
x"00",x"00",x"00",x"FD",x"DD",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FD",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FD",x"DC",x"DC",x"DC",x"FD",x"00",x"00",
x"00",x"00",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"FD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DD",x"DC",x"FD",x"FE",x"DD",x"DD",x"DD",x"00",
x"00",x"FE",x"DD",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"DD",x"DC",x"FD",x"00",
x"00",x"00",x"FE",x"DC",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"00",x"DC",x"DD",x"00",x"FE",
x"DC",x"DD",x"00",x"00",x"DC",x"FD",x"00",x"DD",
x"DC",x"DD",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FD",x"DC",x"DD",x"DD",x"FE",x"00",x"00",x"00",
x"00",x"DD",x"FE",x"DD",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"DD",x"DC",x"FE",x"00",x"00",
x"00",x"00",x"DD",x"DC",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"FE",
x"DD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"FE",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"DD",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DD",x"DC",x"00",x"00",x"00",
x"FE",x"DD",x"DC",x"FE",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"FD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"DD",x"DC",x"DC",x"DC",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",
x"00",x"00",x"DD",x"DC",x"00",x"00",x"00",x"00",
x"FE",x"DD",x"00",x"00",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"FD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FE",x"FE",x"FE",x"FE",x"FD",x"DD",x"DC",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",
x"00",x"FE",x"DC",x"DC",x"00",x"00",x"00",x"FE",
x"DC",x"DD",x"FE",x"FE",x"DC",x"DD",x"FE",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"FE",
x"DD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"FE",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DD",x"FE",x"DD",x"DD",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"00",
x"DD",x"DD",x"DD",x"DD",x"DC",x"DC",x"FE",x"00",
x"00",x"00",x"00",x"00",x"DC",x"DD",x"00",x"FE",
x"DC",x"DD",x"00",x"00",x"DC",x"FD",x"00",x"DD",
x"DC",x"DD",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FD",x"DC",x"DC",x"DC",x"FD",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",
x"00",x"FE",x"DC",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"DC",x"DD",x"00",x"FE",
x"DC",x"DC",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"FD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FD",x"FE",x"00",x"00",x"00",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
); 


  constant ROM_CAR : type_ROM := 
(x"DC",x"94",x"00",x"00",x"24",x"B4",x"DC",x"B8",
x"00",x"00",x"6C",x"DC",x"DC",x"04",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D8",x"DC",x"90",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"90",x"DC",x"DC",
x"DC",x"B8",x"48",x"00",x"90",x"DC",x"DC",x"B8",
x"00",x"00",x"6C",x"DC",x"70",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D8",x"DC",x"90",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"90",x"DC",x"DC",
x"B8",x"DC",x"90",x"00",x"90",x"DC",x"B8",x"B8",
x"00",x"00",x"6C",x"DC",x"24",x"00",x"24",x"B8",
x"B8",x"B8",x"4C",x"00",x"00",x"D8",x"DC",x"90",
x"00",x"00",x"90",x"B8",x"B8",x"B8",x"90",x"00",
x"00",x"00",x"94",x"B8",x"B8",x"B8",x"6C",x"00",
x"00",x"90",x"B8",x"B8",x"B8",x"B8",x"B8",x"48",
x"90",x"B8",x"B8",x"90",x"00",x"00",x"00",x"90",
x"B8",x"B8",x"90",x"00",x"00",x"90",x"DC",x"DC",
x"00",x"DC",x"90",x"24",x"B4",x"DC",x"00",x"DC",
x"B4",x"48",x"DC",x"DC",x"24",x"48",x"DC",x"B8",
x"70",x"B4",x"DC",x"70",x"00",x"D8",x"DC",x"90",
x"00",x"70",x"DC",x"90",x"70",x"DC",x"DC",x"70",
x"00",x"90",x"DC",x"70",x"70",x"94",x"DC",x"90",
x"04",x"B4",x"DC",x"D8",x"70",x"94",x"DC",x"DC",
x"90",x"70",x"DC",x"B8",x"24",x"24",x"B4",x"DC",
x"90",x"90",x"DC",x"B4",x"24",x"48",x"B8",x"DC",
x"00",x"DC",x"90",x"6C",x"DC",x"6C",x"00",x"DC",
x"B4",x"48",x"DC",x"70",x"00",x"B8",x"DC",x"D8",
x"94",x"B8",x"DC",x"DC",x"24",x"D8",x"DC",x"90",
x"48",x"B8",x"DC",x"24",x"00",x"28",x"28",x"24",
x"48",x"D8",x"DC",x"00",x"00",x"00",x"70",x"DC",
x"48",x"B4",x"DC",x"B4",x"00",x"48",x"DC",x"DC",
x"24",x"00",x"DC",x"DC",x"90",x"6C",x"DC",x"DC",
x"94",x"94",x"DC",x"DC",x"6C",x"00",x"B4",x"48",
x"00",x"DC",x"DC",x"DC",x"DC",x"24",x"00",x"94",
x"DC",x"DC",x"DC",x"48",x"00",x"B8",x"DC",x"D8",
x"94",x"94",x"94",x"94",x"00",x"D8",x"DC",x"90",
x"4C",x"DC",x"DC",x"24",x"00",x"00",x"00",x"00",
x"70",x"DC",x"DC",x"00",x"00",x"00",x"4C",x"DC",
x"48",x"B4",x"DC",x"B4",x"00",x"48",x"DC",x"DC",
x"24",x"00",x"DC",x"DC",x"90",x"6C",x"DC",x"DC",
x"94",x"94",x"94",x"94",x"48",x"00",x"94",x"00",
x"00",x"70",x"DC",x"DC",x"DC",x"24",x"00",x"00",
x"DC",x"DC",x"DC",x"48",x"00",x"B8",x"DC",x"B4",
x"00",x"24",x"70",x"70",x"00",x"D8",x"DC",x"90",
x"24",x"B4",x"DC",x"24",x"00",x"00",x"70",x"48",
x"24",x"B4",x"DC",x"00",x"00",x"24",x"94",x"DC",
x"48",x"B4",x"DC",x"B4",x"00",x"48",x"DC",x"DC",
x"24",x"00",x"DC",x"DC",x"90",x"6C",x"DC",x"DC",
x"00",x"00",x"70",x"70",x"28",x"00",x"48",x"00",
x"00",x"24",x"DC",x"DC",x"6C",x"00",x"00",x"00",
x"DC",x"DC",x"70",x"00",x"00",x"00",x"B8",x"D8",
x"B8",x"D8",x"D8",x"48",x"00",x"D8",x"DC",x"90",
x"00",x"6C",x"D8",x"B8",x"B8",x"B8",x"D8",x"6C",
x"00",x"70",x"D8",x"B8",x"B8",x"B8",x"D8",x"6C",
x"00",x"B4",x"DC",x"B4",x"00",x"48",x"DC",x"DC",
x"24",x"00",x"DC",x"DC",x"90",x"00",x"90",x"D8",
x"B8",x"B8",x"D8",x"70",x"00",x"6C",x"B8",x"B8",
x"00",x"04",x"70",x"70",x"24",x"00",x"00",x"00",
x"70",x"70",x"28",x"00",x"00",x"00",x"00",x"70",
x"70",x"70",x"24",x"00",x"00",x"6C",x"70",x"48",
x"00",x"00",x"48",x"70",x"70",x"70",x"48",x"00",
x"00",x"00",x"6C",x"70",x"70",x"70",x"48",x"00",
x"00",x"6C",x"70",x"6C",x"00",x"24",x"70",x"70",
x"00",x"00",x"70",x"70",x"48",x"00",x"00",x"4C",
x"70",x"70",x"4C",x"00",x"00",x"48",x"70",x"70",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"24",x"4C",x"4C",x"4C",x"4C",x"48",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"24",x"B4",x"DC",x"DC",x"DC",x"DC",x"D8",
x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"B8",x"48",x"00",x"00",x"90",x"DC",
x"D8",x"6C",x"00",x"00",x"24",x"28",x"28",x"28",
x"24",x"00",x"00",x"24",x"28",x"28",x"28",x"24",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"90",x"DC",x"90",x"00",x"00",x"00",x"00",x"4C",
x"48",x"00",x"00",x"48",x"B8",x"DC",x"DC",x"DC",
x"90",x"00",x"00",x"94",x"DC",x"DC",x"DC",x"90",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DC",x"DC",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"6C",x"B8",x"48",x"48",x"DC",
x"D8",x"6C",x"00",x"94",x"DC",x"24",x"04",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DC",x"DC",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"24",x"4C",x"D8",x"DC",x"DC",
x"DC",x"6C",x"00",x"94",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"48",x"DC",x"90",x"00",x"00",x"00",x"00",x"94",
x"6C",x"00",x"48",x"B8",x"DC",x"48",x"48",x"DC",
x"DC",x"6C",x"00",x"94",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"B4",x"DC",x"90",x"28",x"28",x"B8",x"DC",
x"D8",x"6C",x"6C",x"DC",x"DC",x"48",x"48",x"DC",
x"DC",x"6C",x"00",x"94",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"90",x"DC",x"DC",x"DC",x"DC",x"D8",
x"48",x"00",x"24",x"B4",x"DC",x"DC",x"D8",x"6C",
x"DC",x"6C",x"00",x"94",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"00",
x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",
x"04",x"00",x"00",x"00",x"04",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"B8",x"B8",x"B8",x"B8",x"B8",x"B8",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B8",
x"B8",x"6C",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"B8",x"70",x"70",x"70",x"D8",x"D8",
x"48",x"00",x"00",x"00",x"00",x"00",x"00",x"70",
x"70",x"48",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"90",x"00",x"00",x"00",x"24",x"DC",
x"B4",x"00",x"48",x"94",x"94",x"94",x"94",x"94",
x"94",x"48",x"00",x"00",x"70",x"94",x"94",x"94",
x"48",x"00",x"00",x"00",x"90",x"94",x"94",x"48",
x"00",x"00",x"00",x"90",x"94",x"6C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"94",x"28",x"28",x"28",x"B8",x"D8",
x"6C",x"00",x"6C",x"DC",x"B4",x"94",x"94",x"DC",
x"DC",x"6C",x"00",x"94",x"DC",x"94",x"B4",x"DC",
x"DC",x"4C",x"24",x"B8",x"DC",x"94",x"B4",x"DC",
x"70",x"00",x"00",x"90",x"94",x"6C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"48",
x"00",x"00",x"6C",x"DC",x"24",x"00",x"00",x"DC",
x"DC",x"6C",x"48",x"B8",x"DC",x"00",x"00",x"4C",
x"4C",x"24",x"90",x"DC",x"D8",x"70",x"94",x"DC",
x"DC",x"48",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"90",x"04",x"04",x"04",x"04",x"00",
x"00",x"00",x"6C",x"DC",x"24",x"00",x"00",x"DC",
x"DC",x"6C",x"70",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"94",x"DC",x"DC",x"B8",x"B8",x"B8",
x"B8",x"24",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"6C",x"DC",x"24",x"00",x"00",x"DC",
x"DC",x"6C",x"48",x"B8",x"DC",x"00",x"00",x"04",
x"4C",x"24",x"90",x"DC",x"D8",x"00",x"00",x"4C",
x"4C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"6C",x"DC",x"24",x"00",x"00",x"DC",
x"DC",x"6C",x"00",x"94",x"DC",x"94",x"94",x"B4",
x"DC",x"4C",x"24",x"B8",x"DC",x"94",x"B4",x"DC",
x"70",x"00",x"00",x"90",x"94",x"6C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"94",x"4C",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"48",x"94",x"24",x"00",x"00",x"94",
x"94",x"48",x"00",x"00",x"70",x"94",x"94",x"94",
x"48",x"00",x"00",x"00",x"90",x"94",x"94",x"48",
x"00",x"00",x"00",x"90",x"94",x"6C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"28",x"90",x"6C",x"00",x"00",x"00",
x"00",x"00",x"00",x"24",x"28",x"00",x"00",x"00",
x"28",x"28",x"28",x"28",x"28",x"28",x"24",x"00",
x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"28",
x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"28",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"90",x"DC",x"DC",x"DC",x"90",x"00",x"00",
x"00",x"00",x"24",x"B4",x"DC",x"04",x"00",x"24",
x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"B4",x"00",
x"00",x"00",x"00",x"6C",x"D8",x"B4",x"00",x"00",
x"00",x"00",x"00",x"00",x"90",x"DC",x"DC",x"DC",
x"94",x"00",x"00",x"00",x"90",x"DC",x"DC",x"DC",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"B8",x"DC",x"90",x"70",x"D8",x"B8",x"94",x"00",
x"00",x"48",x"D8",x"DC",x"DC",x"04",x"00",x"00",
x"04",x"04",x"04",x"24",x"B8",x"DC",x"90",x"00",
x"00",x"00",x"70",x"D8",x"DC",x"B4",x"00",x"00",
x"00",x"00",x"00",x"24",x"DC",x"94",x"04",x"90",
x"DC",x"B8",x"00",x"24",x"DC",x"90",x"04",x"94",
x"DC",x"B8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"90",x"DC",x"B4",x"94",x"48",x"00",x"00",x"00",
x"24",x"B8",x"70",x"B4",x"DC",x"04",x"00",x"00",
x"00",x"00",x"00",x"94",x"DC",x"6C",x"00",x"00",
x"00",x"24",x"B4",x"DC",x"DC",x"B4",x"00",x"00",
x"00",x"00",x"00",x"D8",x"DC",x"90",x"00",x"48",
x"B8",x"DC",x"00",x"DC",x"DC",x"70",x"00",x"48",
x"B8",x"D8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"B4",x"24",x"00",x"00",
x"00",x"24",x"00",x"90",x"DC",x"04",x"00",x"00",
x"00",x"00",x"48",x"D8",x"DC",x"00",x"00",x"00",
x"48",x"B8",x"DC",x"48",x"D8",x"B4",x"00",x"00",
x"00",x"00",x"00",x"D8",x"DC",x"90",x"00",x"00",
x"90",x"DC",x"00",x"DC",x"DC",x"70",x"00",x"00",
x"B4",x"D8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"24",x"B8",x"DC",x"DC",x"DC",x"00",
x"00",x"00",x"00",x"90",x"DC",x"04",x"00",x"00",
x"00",x"00",x"94",x"DC",x"24",x"00",x"00",x"00",
x"90",x"B4",x"24",x"00",x"D8",x"B4",x"00",x"00",
x"00",x"00",x"00",x"D8",x"DC",x"90",x"00",x"00",
x"90",x"DC",x"00",x"DC",x"DC",x"70",x"00",x"00",
x"B4",x"D8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"70",x"70",x"48",x"6C",x"90",x"B8",x"DC",x"00",
x"00",x"00",x"00",x"90",x"DC",x"04",x"00",x"00",
x"00",x"6C",x"DC",x"DC",x"24",x"00",x"00",x"48",
x"DC",x"94",x"70",x"70",x"D8",x"D8",x"48",x"00",
x"00",x"00",x"00",x"D8",x"DC",x"90",x"00",x"48",
x"B8",x"DC",x"00",x"DC",x"DC",x"70",x"00",x"48",
x"B8",x"D8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"24",x"DC",x"D8",x"D8",x"6C",x"B4",x"B8",x"00",
x"00",x"00",x"00",x"90",x"DC",x"04",x"00",x"00",
x"00",x"6C",x"DC",x"48",x"00",x"00",x"00",x"28",
x"B8",x"B8",x"B8",x"B8",x"DC",x"D8",x"70",x"00",
x"04",x"04",x"00",x"24",x"DC",x"94",x"04",x"90",
x"DC",x"B8",x"00",x"28",x"DC",x"90",x"04",x"94",
x"DC",x"B8",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"90",x"DC",x"DC",x"DC",x"90",x"00",x"00",
x"00",x"00",x"00",x"90",x"DC",x"04",x"00",x"00",
x"00",x"6C",x"DC",x"28",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D8",x"B4",x"00",x"4C",
x"DC",x"DC",x"24",x"00",x"90",x"DC",x"DC",x"DC",
x"94",x"00",x"00",x"00",x"90",x"DC",x"DC",x"DC",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"28",x"90",x"70",x"00",x"00",x"00",
x"48",x"00",x"00",x"24",x"28",x"00",x"00",x"00",
x"00",x"00",x"28",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",
x"28",x"28",x"00",x"00",x"00",x"28",x"28",x"28",
x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"28",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
); 


  constant ROM_TRUCK : type_ROM := 
(x"DC",x"DD",x"00",x"00",x"00",x"DD",x"DC",x"DD",
x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FD",x"DC",x"DC",
x"DC",x"DD",x"FE",x"00",x"FD",x"DC",x"DC",x"DD",
x"00",x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FD",x"DC",x"DC",
x"DD",x"DC",x"FD",x"00",x"FD",x"DC",x"DD",x"DD",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DD",
x"DD",x"DD",x"FE",x"00",x"00",x"DC",x"DC",x"FD",
x"00",x"00",x"FE",x"DD",x"DD",x"DD",x"FE",x"00",
x"00",x"00",x"FD",x"DD",x"DD",x"DD",x"FE",x"00",
x"00",x"FD",x"DD",x"DD",x"DD",x"DD",x"DD",x"FE",
x"FD",x"DD",x"DD",x"FE",x"00",x"00",x"00",x"FD",
x"DD",x"DD",x"FD",x"00",x"00",x"FD",x"DC",x"DC",
x"00",x"DC",x"FD",x"00",x"DD",x"DC",x"00",x"DC",
x"DD",x"FE",x"DC",x"DC",x"00",x"00",x"DC",x"DD",
x"FD",x"DD",x"DC",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"FE",x"DC",x"DD",x"FD",x"DC",x"DC",x"FE",
x"00",x"FD",x"DC",x"FD",x"FD",x"DD",x"DC",x"FD",
x"00",x"DD",x"DC",x"DC",x"FD",x"DD",x"DC",x"DC",
x"DD",x"FD",x"DC",x"DD",x"00",x"00",x"DD",x"DC",
x"FD",x"FD",x"DC",x"DD",x"00",x"FE",x"DD",x"DC",
x"00",x"DC",x"FD",x"FE",x"DC",x"FE",x"00",x"DC",
x"DD",x"FE",x"DC",x"FD",x"00",x"DD",x"DC",x"DD",
x"FD",x"DD",x"DC",x"DC",x"00",x"DC",x"DC",x"FD",
x"00",x"DD",x"DC",x"00",x"00",x"FE",x"FE",x"00",
x"FE",x"DD",x"DC",x"00",x"00",x"00",x"FD",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"FD",x"FD",x"DC",x"DC",x"FE",x"00",x"DD",x"FE",
x"00",x"DC",x"DC",x"DC",x"DC",x"00",x"00",x"DD",
x"DC",x"DC",x"DC",x"FE",x"00",x"DD",x"DC",x"DC",
x"DD",x"DD",x"DD",x"DD",x"00",x"DC",x"DC",x"FD",
x"FE",x"DC",x"DC",x"00",x"00",x"00",x"00",x"00",
x"FE",x"DC",x"DC",x"00",x"00",x"00",x"FE",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"DD",x"DD",x"DD",x"DD",x"FE",x"00",x"DD",x"00",
x"00",x"FD",x"DC",x"DC",x"DC",x"00",x"00",x"00",
x"DC",x"DC",x"DC",x"FE",x"00",x"DD",x"DC",x"DD",
x"00",x"00",x"FE",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"DD",x"DC",x"00",x"00",x"00",x"FE",x"00",
x"FE",x"DD",x"DC",x"00",x"00",x"00",x"FD",x"DC",
x"FE",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"FE",x"DC",x"DC",
x"00",x"00",x"FE",x"FE",x"00",x"00",x"FE",x"00",
x"00",x"00",x"DC",x"DC",x"FE",x"00",x"00",x"00",
x"DC",x"DC",x"FD",x"00",x"00",x"00",x"DC",x"DC",
x"DD",x"DD",x"DC",x"FE",x"00",x"DC",x"DC",x"FD",
x"00",x"FE",x"DC",x"DD",x"DD",x"DD",x"DC",x"FE",
x"00",x"FD",x"DC",x"DD",x"DD",x"DD",x"DC",x"FE",
x"00",x"DD",x"DC",x"DD",x"00",x"FE",x"DC",x"DC",
x"00",x"00",x"DC",x"DC",x"FE",x"00",x"DD",x"DC",
x"DD",x"DD",x"DC",x"DD",x"00",x"FE",x"DD",x"DD",
x"00",x"00",x"DD",x"DD",x"00",x"00",x"00",x"00",
x"DD",x"DD",x"FE",x"00",x"00",x"00",x"00",x"DD",
x"DD",x"DD",x"FE",x"00",x"00",x"DD",x"DD",x"FE",
x"00",x"00",x"FE",x"DD",x"DD",x"DD",x"FE",x"00",
x"00",x"00",x"FE",x"DD",x"DD",x"DD",x"FE",x"00",
x"00",x"FE",x"DD",x"FD",x"00",x"00",x"DD",x"DD",
x"00",x"00",x"DD",x"DD",x"FE",x"00",x"00",x"FE",
x"DD",x"DD",x"FE",x"00",x"00",x"FE",x"DD",x"DD",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FD",x"DC",x"DC",x"FE",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"DC",x"DC",x"DC",x"00",x"DC",
x"FD",x"00",x"00",x"FD",x"DC",x"DD",x"00",x"00",
x"FE",x"DC",x"DC",x"DC",x"DD",x"00",x"00",x"FE",
x"DC",x"FE",x"00",x"DD",x"DC",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"FD",x"FE",x"FE",x"00",x"DC",
x"FD",x"00",x"00",x"DD",x"DC",x"DD",x"00",x"FE",
x"DC",x"DD",x"FE",x"DD",x"DC",x"DD",x"00",x"FE",
x"DC",x"FD",x"DD",x"DC",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"DC",
x"FD",x"00",x"00",x"DD",x"DC",x"DD",x"00",x"DD",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"FE",
x"DC",x"DC",x"DC",x"DC",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"DC",
x"FD",x"00",x"00",x"DD",x"DC",x"DD",x"00",x"DC",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"FE",
x"DC",x"DC",x"DC",x"DC",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"DC",
x"FD",x"00",x"00",x"DD",x"DC",x"DD",x"00",x"FE",
x"DC",x"FE",x"00",x"00",x"FE",x"FE",x"00",x"FE",
x"DC",x"FE",x"FE",x"DC",x"DD",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DC",x"DC",x"00",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"DD",
x"DC",x"DD",x"DD",x"DC",x"DC",x"DD",x"00",x"00",
x"DD",x"DD",x"DD",x"DD",x"DC",x"FD",x"00",x"FE",
x"DC",x"FE",x"00",x"DD",x"DC",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FE",x"FD",x"00",x"00",
x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"00",
x"00",x"FE",x"FE",x"FE",x"FE",x"00",x"00",x"00",
x"FE",x"00",x"00",x"00",x"FE",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"FE",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"DD",x"DC",
x"FD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"FE",x"DC",
x"DD",x"00",x"FE",x"DC",x"DC",x"DC",x"DC",x"DC",
x"DC",x"FE",x"00",x"00",x"DD",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"FE",x"DC",x"DC",x"DC",x"DD",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DD",x"FD",x"FD",x"FD",x"DC",x"DD",
x"00",x"00",x"FE",x"DC",x"FE",x"FE",x"FE",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"FE",x"FE",x"DC",
x"DC",x"FE",x"FE",x"DC",x"DC",x"FE",x"FE",x"DC",
x"DD",x"00",x"00",x"FE",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DD",x"DD",x"DD",x"DD",x"DD",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"FE",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"FD",x"DC",x"DC",x"DC",x"DC",x"DC",
x"DC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"FE",x"DC",x"DC",x"00",x"00",x"00",
x"00",x"00",x"FD",x"DC",x"DC",x"FE",x"FE",x"FE",
x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"00",x"DD",x"DC",x"00",x"00",x"00",
x"DD",x"FE",x"FD",x"DC",x"DC",x"00",x"00",x"DD",
x"DD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"FD",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"00",x"00",x"00",x"DC",
x"DC",x"FE",x"00",x"FE",x"DC",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"FE",x"DC",x"DC",x"DC",x"DD",
x"FE",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"FE",
x"FE",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"FE",
x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"00",
x"00",x"00",x"00",x"FE",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DD",x"FD",x"00",x"00",x"00",
x"00",x"00",x"FE",x"FE",x"FE",x"00",x"00",x"00",
x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",
x"00",x"00",x"FE",x"FE",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",
x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"DC",x"DC",x"DC",x"DD",x"00",x"00",
x"00",x"DD",x"DC",x"DC",x"DC",x"DD",x"00",x"00",
x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"00",
x"FE",x"DD",x"DC",x"DC",x"DC",x"FE",x"00",x"00",
x"00",x"00",x"00",x"00",x"DD",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"00",x"DD",x"DC",x"DC",x"DC",
x"DD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"DC",x"DC",x"FD",x"FE",x"DD",x"DD",x"DD",x"00",
x"00",x"DD",x"FE",x"00",x"DD",x"DC",x"00",x"00",
x"00",x"00",x"00",x"00",x"DD",x"DC",x"FE",x"00",
x"FE",x"DC",x"00",x"00",x"DC",x"DC",x"FD",x"00",
x"00",x"00",x"00",x"00",x"DC",x"FD",x"00",x"FE",
x"DC",x"DC",x"00",x"FE",x"DC",x"FE",x"00",x"FD",
x"DC",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FE",x"DC",x"DD",x"DD",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"DD",x"DC",x"00",x"00",
x"00",x"00",x"00",x"DD",x"DC",x"FE",x"00",x"00",
x"FE",x"DC",x"00",x"00",x"DC",x"DC",x"FD",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"DD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"DC",x"DC",x"DD",x"00",x"00",x"00",
x"00",x"00",x"FE",x"DD",x"DC",x"DC",x"00",x"00",
x"00",x"00",x"FE",x"DC",x"DD",x"00",x"00",x"00",
x"00",x"FD",x"DD",x"DD",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"FD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"DD",x"DC",x"DC",x"DC",x"00",
x"00",x"00",x"00",x"00",x"FE",x"DC",x"DD",x"00",
x"00",x"00",x"DD",x"DC",x"00",x"00",x"00",x"00",
x"FE",x"DC",x"DD",x"FD",x"DC",x"DD",x"00",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"00",
x"FD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FD",x"FD",x"FE",x"FE",x"FE",x"DD",x"DC",x"00",
x"FD",x"FD",x"FE",x"00",x"00",x"DD",x"DD",x"00",
x"00",x"FE",x"DC",x"DC",x"00",x"00",x"00",x"00",
x"DD",x"DC",x"00",x"00",x"FE",x"DC",x"FD",x"00",
x"00",x"00",x"00",x"DC",x"DC",x"FD",x"00",x"FE",
x"DD",x"DC",x"00",x"DC",x"DC",x"FE",x"00",x"FE",
x"DD",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"DC",x"DC",x"DC",x"FE",x"DD",x"DD",x"00",
x"DD",x"DC",x"FE",x"00",x"DD",x"DC",x"DD",x"00",
x"00",x"FE",x"DC",x"FE",x"00",x"00",x"00",x"00",
x"DD",x"DC",x"FE",x"00",x"DD",x"DC",x"FE",x"00",
x"00",x"00",x"00",x"00",x"DC",x"DD",x"00",x"FD",
x"DC",x"DD",x"00",x"00",x"DC",x"FD",x"00",x"DD",
x"DC",x"DD",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FD",x"DC",x"DC",x"DC",x"FD",x"00",x"00",
x"00",x"DD",x"DC",x"DC",x"DC",x"FE",x"00",x"00",
x"00",x"FE",x"DC",x"00",x"00",x"00",x"00",x"00",
x"00",x"DD",x"DC",x"DC",x"DC",x"FE",x"00",x"FE",
x"DC",x"DC",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"FD",x"00",x"00",x"00",x"FD",x"DC",x"DC",x"DC",
x"FD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FD",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
); 

  constant ROM_GO : type_ROM := 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",
x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"48",x"6C",x"90",x"B4",x"B4",
x"B4",x"B4",x"90",x"48",x"24",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"6C",x"90",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"48",x"90",x"94",x"B4",x"90",x"90",
x"90",x"90",x"B4",x"94",x"6C",x"24",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"90",x"D9",
x"B9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"24",x"B4",x"D9",x"90",x"48",x"00",x"00",
x"00",x"24",x"6C",x"B9",x"B4",x"6C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"90",x"D9",
x"B9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"28",x"90",x"DD",x"48",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"6C",x"B4",x"D9",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"90",x"D9",
x"B9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"6C",x"B4",x"B5",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"24",x"48",x"6C",x"00",x"00",
x"00",x"00",x"48",x"90",x"B4",x"B5",x"B5",x"B4",
x"90",x"24",x"00",x"00",x"00",x"00",x"90",x"B9",
x"B4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"90",x"B9",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",
x"00",x"24",x"94",x"B4",x"94",x"70",x"70",x"94",
x"B4",x"90",x"24",x"00",x"00",x"00",x"90",x"B5",
x"B4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"94",x"B9",x"6C",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"04",x"6C",x"D9",x"90",x"48",x"00",x"00",x"48",
x"90",x"DD",x"48",x"04",x"00",x"00",x"70",x"B4",
x"94",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",
x"94",x"B5",x"48",x"00",x"00",x"00",x"00",x"00",
x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",
x"24",x"B5",x"94",x"28",x"00",x"00",x"00",x"00",
x"24",x"D9",x"90",x"48",x"00",x"00",x"6C",x"94",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",
x"94",x"B9",x"48",x"00",x"00",x"00",x"00",x"48",
x"90",x"D9",x"D9",x"D9",x"D9",x"B9",x"48",x"00",
x"48",x"D9",x"6C",x"24",x"00",x"00",x"00",x"00",
x"00",x"94",x"B4",x"4C",x"00",x"00",x"6C",x"90",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"90",x"B9",x"6C",x"00",x"00",x"00",x"00",x"24",
x"48",x"6C",x"6C",x"6C",x"94",x"DD",x"4C",x"24",
x"48",x"DD",x"4C",x"24",x"00",x"00",x"00",x"00",
x"00",x"90",x"B4",x"6C",x"00",x"00",x"6C",x"90",
x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"90",x"B9",x"90",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"6C",x"DD",x"4C",x"24",
x"48",x"DD",x"6C",x"24",x"00",x"00",x"00",x"00",
x"00",x"90",x"B4",x"6C",x"00",x"00",x"48",x"6C",
x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"6C",x"B4",x"D9",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"6C",x"DD",x"4C",x"04",
x"48",x"D9",x"70",x"24",x"00",x"00",x"00",x"00",
x"00",x"B4",x"94",x"48",x"00",x"00",x"24",x"48",
x"48",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"04",x"4C",x"DD",x"94",x"48",x"00",x"00",x"00",
x"00",x"00",x"00",x"48",x"90",x"DD",x"4C",x"00",
x"24",x"90",x"B9",x"48",x"00",x"00",x"00",x"00",
x"48",x"DD",x"70",x"24",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"24",x"6C",x"B5",x"94",x"70",x"48",x"48",
x"48",x"48",x"70",x"94",x"B4",x"B4",x"24",x"00",
x"00",x"48",x"D9",x"94",x"6C",x"48",x"48",x"6C",
x"94",x"B9",x"48",x"00",x"00",x"00",x"48",x"6C",
x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"24",x"90",x"94",x"B4",x"90",x"90",
x"90",x"90",x"B4",x"B4",x"90",x"4C",x"00",x"00",
x"00",x"00",x"90",x"94",x"B4",x"90",x"90",x"94",
x"B4",x"6C",x"00",x"00",x"00",x"00",x"70",x"B4",
x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"24",x"6C",x"90",x"B4",
x"B4",x"94",x"6C",x"24",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"48",x"70",x"B4",x"94",x"70",
x"48",x"00",x"00",x"00",x"00",x"00",x"48",x"4C",
x"48",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
); 

  signal Location : natural range 0 to 65535;  

begin
	  
  --Address <= Xin(5 downto 0) + (Yin(5 downto 0)&"000000");
  --Address <= (conv_integer(Xin(5 downto 0))) - 288 + (conv_integer(Yin(5 downto 0)&"000000")-208);
  Address <= (conv_integer(Xin) - 288) + (conv_integer((Yin(5 downto 0)-208)&"000000"));

  process (Clk)
  begin
    -- Check if pixel is in the active zone
	 if rising_edge(Clk) then
	   if (En = '1') then
	     if ((Xin>=288 and Xin < 352) and (Yin>=208 and Yin < 272)) then
			    case (img) is 
					when "000" =>
						Color <= ROM_MOTORCYCLE (Address);
					when "001" =>
						Color <= ROM_CAR (Address);
					when "010" =>
						Color <= ROM_CAR (Address);
					when "011" =>
						Color <= ROM_TRUCK (Address);
					when "100" =>
						Color <= ROM_GO (Address);
					when others =>
						Color <= ROM_MOTORCYCLE (Address);
					end case;
		  else
          Color <= "00000000"; -- Black
		  end if;
		else 
		  Color <= "00000000"; -- Black
	   end if;
	 end if;
  end process;
  
  -- Send individual color to their channel
  R <= Color(7 downto 5);
  G <= Color(4 downto 2);
  B <= Color(1 downto 0);

end Behavioral;


